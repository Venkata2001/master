// Code your testbench here
// or browse Examples
`include "i3c_top.sv"
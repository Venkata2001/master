typedef uvm_sequencer#(base_tx) s_seq;
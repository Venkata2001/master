class base_tx extends uvm_sequence_item;
`uvm_object_utils(base_tx)
`NEW_OBJ
endclass

class env_cfg extends uvm_object;
  `uvm_object_utils(env_cfg)
  `NEW_OBJ
  //seting no_of_slaves
  int no_of_slaves=5; 
endclass
typedef uvm_sequencer#(base_tx) m_seq;
